/nethome/mi72/sideProjects/Fibonacci-Circuit/src/uvm/sequences/fibonacci_seq_lib.sv