/nethome/mi72/sideProjects/Fibonacci-Circuit/src/uvm/tests/fibonacci_test_lib.sv