package fibonacci_seq_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "fibonacci_seq_item.sv"
  `include "fibonacci_sequence.svh"
  `include "fibonacci_seq_lib.sv"
  
endpackage : fibonacci_seq_pkg
