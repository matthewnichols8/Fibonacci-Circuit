/nethome/mi72/sideProjects/Fibonacci-Circuit/src/uvm/agent/fibonacci_agent.sv