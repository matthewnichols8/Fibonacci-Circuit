package fibonacci_test_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import fibonacci_env_pkg::*;
  import fibonacci_seq_pkg::*;
  `include "fibonacci_base_test.svh"
  `include "fibonacci_test_lib.sv"
  
endpackage : fibonacci_test_pkg
