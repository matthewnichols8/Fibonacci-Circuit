/nethome/mi72/sideProjects/Fibonacci-Circuit/src/uvm/tb/fibonacci_if.sv