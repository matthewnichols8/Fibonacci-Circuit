/nethome/mi72/sideProjects/Fibonacci-Circuit/src/uvm/env/fibonacci_env.sv