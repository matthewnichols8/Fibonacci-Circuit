/nethome/mi72/sideProjects/Fibonacci-Circuit/src/sv/rtl/fibonacci.sv