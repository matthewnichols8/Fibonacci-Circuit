/nethome/mi72/sideProjects/Fibonacci-Circuit/src/uvm/tests/fibonacci_base_test.svh